`timescale 1ns/1ns
module SixteenBarrelShifter(input [15:0] A,input [3:0] N,output [15:0] w);
	SixteenMux CUT1({A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14]},N,w[15]);
	SixteenMux CUT2({A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13]},N,w[14]);
	SixteenMux CUT3({A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12]},N,w[13]);
	SixteenMux CUT4({A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11]},N,w[12]);
	SixteenMux CUT5({A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10]},N,w[11]);
	SixteenMux CUT6({A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9]},N,w[10]);
	SixteenMux CUT7({A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8]},N,w[9]);
	SixteenMux CUT8({A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7]},N,w[8]);
	SixteenMux CUT9({A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5],A[6]},N,w[7]);
	SixteenMux CUT10({A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4],A[5]},N,w[6]);
	SixteenMux CUT11({A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3],A[4]},N,w[5]);
	SixteenMux CUT12({A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2],A[3]},N,w[4]);
	SixteenMux CUT13({A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1],A[2]},N,w[3]);
	SixteenMux CUT14({A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0],A[1]},N,w[2]);
	SixteenMux CUT15({A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15],A[0]},N,w[1]);
	SixteenMux CUT16({A[0],A[1],A[2],A[3],A[4],A[5],A[6],A[7],A[8],A[9],A[10],A[11],A[12],A[13],A[14],A[15]},N,w[0]);
endmodule