`timescale 1ns/1ns
module MUXComparison();
	wire mux1_output,mux2_output;
	reg ss0,ss1,aa,bb,cc,dd;
	MyMUX mux1(ss0,ss1,aa,bb,cc,dd,mux1_output);
	MyMUX2 mux2(ss0,ss1,aa,bb,cc,dd,mux2_output);
	initial begin
	#10 ss0 = 1;ss1 = 1; aa = 0;bb = 0; cc = 0;dd = 1;
	#30
	#15 ss0 = 1;ss1 = 0; aa = 1;bb = 0; cc = 0;dd = 1;
	#20
	#30 $stop;
	end
endmodule